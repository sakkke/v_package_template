module v_package_template

fn hello() {
	println('Hello World!')
}
